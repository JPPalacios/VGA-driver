--> in-progress

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

package vga_pkg is





end package;

package body vga_pkg is

end package body;